----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/31/2025 12:48:12 PM
-- Design Name: 
-- Module Name: riconoscitore_101 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity riconoscitore_101 is
    Port (  input   :   in  std_logic;
            a       :   in  std_logic; -- segnale ti tempificazione(clock)
            reset   :   in  std_logic;
            m       :   in  std_logic; --0 modalità non sovrapposta, 1 modalità parzialmente sovrapposta
            output  :   out std_logic
     );
end riconoscitore_101;

architecture Behavioral of riconoscitore_101 is
    
    type    stato is (S0,S1,S2);
    signal  stato_corrente  :   stato   :=S0;
    signal  stato_prossimo  :   stato;
begin
    
    state_proccess: process(stato_corrente,input,m)
        begin
            if(m)   then 
                case stato_corrente is
                    when    
                end case;
            else
                case stato_corrente is
                    when    
                end case;
    end process;
    
    memory_process  :   process (a)
        begin   
            if(a'event and a='1')   then
                stato_corrente<=stato_prossimo;
            end if;
    end process;


end Behavioral;
